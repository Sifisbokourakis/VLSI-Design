** Profile: "SCHEMATIC1-DC"  [ C:\Users\VLSI_A\Documents\ORCAD\DESIGNS\VLSI-21\Test-PSpiceFiles\SCHEMATIC1\DC.sim ] 

** Creating circuit file "DC.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Cadence/SPB_16.5/tools/pspice/library/UMC_018-TT.lib" 
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V2 0 1.8 10m 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
