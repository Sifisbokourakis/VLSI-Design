** Profile: "VERIFY-Time"  [ C:\Cadence\Designs\VLSI-21\VLSI-21\datapath-pspicefiles\verify\time.sim ] 

** Creating circuit file "Time.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "C:\Cadence\SPB_16.5\tools\pspice\library\UMC 180nm.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 8ns 0 1p 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\VERIFY.net" 


.END
